library verilog;
use verilog.vl_types.all;
entity questao01Arq_vlg_vec_tst is
end questao01Arq_vlg_vec_tst;
