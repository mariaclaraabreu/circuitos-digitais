library verilog;
use verilog.vl_types.all;
entity questao05Arq_vlg_vec_tst is
end questao05Arq_vlg_vec_tst;
