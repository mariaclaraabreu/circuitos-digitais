library verilog;
use verilog.vl_types.all;
entity questao03itema_vlg_check_tst is
    port(
        saida           : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end questao03itema_vlg_check_tst;
