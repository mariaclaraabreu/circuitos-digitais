library verilog;
use verilog.vl_types.all;
entity questao03itemb_vlg_vec_tst is
end questao03itemb_vlg_vec_tst;
