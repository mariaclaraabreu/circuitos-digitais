library verilog;
use verilog.vl_types.all;
entity questao02 is
    port(
        a               : in     vl_logic;
        cicloclk        : in     vl_logic;
        b               : out    vl_logic
    );
end questao02;
