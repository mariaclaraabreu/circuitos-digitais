library verilog;
use verilog.vl_types.all;
entity questao02_vlg_vec_tst is
end questao02_vlg_vec_tst;
