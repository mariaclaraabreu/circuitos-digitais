library verilog;
use verilog.vl_types.all;
entity questao01_vlg_vec_tst is
end questao01_vlg_vec_tst;
