library verilog;
use verilog.vl_types.all;
entity questao04Arq_vlg_check_tst is
    port(
        Saida           : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end questao04Arq_vlg_check_tst;
