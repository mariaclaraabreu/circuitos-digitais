library verilog;
use verilog.vl_types.all;
entity questao04Arq_vlg_vec_tst is
end questao04Arq_vlg_vec_tst;
