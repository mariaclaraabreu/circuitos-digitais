library verilog;
use verilog.vl_types.all;
entity questao03itema_vlg_vec_tst is
end questao03itema_vlg_vec_tst;
