library verilog;
use verilog.vl_types.all;
entity questao01Arq is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        s               : out    vl_logic
    );
end questao01Arq;
