library verilog;
use verilog.vl_types.all;
entity questao02Arq_vlg_vec_tst is
end questao02Arq_vlg_vec_tst;
