library verilog;
use verilog.vl_types.all;
entity questao03Arq_vlg_vec_tst is
end questao03Arq_vlg_vec_tst;
