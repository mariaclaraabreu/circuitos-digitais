library verilog;
use verilog.vl_types.all;
entity questao03Arq is
    port(
        D0              : in     vl_logic;
        D1              : in     vl_logic;
        Sinal           : in     vl_logic;
        Saida           : out    vl_logic
    );
end questao03Arq;
