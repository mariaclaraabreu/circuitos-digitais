library verilog;
use verilog.vl_types.all;
entity questao02Arq_vlg_check_tst is
    port(
        z               : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end questao02Arq_vlg_check_tst;
