library verilog;
use verilog.vl_types.all;
entity questao03itemc_vlg_vec_tst is
end questao03itemc_vlg_vec_tst;
