library verilog;
use verilog.vl_types.all;
entity questao03Arq_vlg_check_tst is
    port(
        Saida           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end questao03Arq_vlg_check_tst;
