library verilog;
use verilog.vl_types.all;
entity questao04Arq_vlg_sample_tst is
    port(
        endereco        : in     vl_logic_vector(2 downto 0);
        sampler_tx      : out    vl_logic
    );
end questao04Arq_vlg_sample_tst;
