library verilog;
use verilog.vl_types.all;
entity questao02_vlg_sample_tst is
    port(
        a               : in     vl_logic;
        cicloclk        : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end questao02_vlg_sample_tst;
