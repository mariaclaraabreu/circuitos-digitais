library verilog;
use verilog.vl_types.all;
entity questao06Arq_vlg_vec_tst is
end questao06Arq_vlg_vec_tst;
